//Verilog HDL for "lab5", "tiehi" "behavioral"


module tiehi_v0( Y );

  output Y;

		assign	Y = 1;


endmodule
