//Verilog HDL for "lab1", "TIELO" "behavioral"
module TIELO ( Y );
  	output Y;
	assign Y = 0;
endmodule
